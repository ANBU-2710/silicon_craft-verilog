module mod_n_count;
endmodule
