module mod_n_count_tb;
endmodule
