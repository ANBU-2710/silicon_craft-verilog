module up_count_tb;
endmodule;
