module down_count;
endmodule
