module up_count;
endmodule
