module piso_tb;
reg clk,rst,shift,load;
reg [width-1:0]
endmodule
