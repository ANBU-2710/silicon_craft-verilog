module down_count_tb;
endmodule
