module ud_count;
endmodule
